typedef uvm_sequencer#(fifo_wtx) fifo_wsqr;
