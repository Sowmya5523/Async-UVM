typedef uvm_sequencer#(fifo_rtx) fifo_rsqr;
